module core;
    initial begin
        $display("Hello, core");
    end
endmodule
