module tb;
    core u_core();
    initial begin
        $display("Hello, World");
        $finish();
    end
endmodule
